`timescale 1ns/1ps

module tb_sha256();
	parameter LOOP = 1;

	reg clk =0;
	//wire [511:0] data = 512'hc13858e5a13de1500e54a1c85f0132e688e131b93d7bf9a00192281e6c555fd0c13858e5a13de1500e54a1c85f0132e688e131b93d7bf9a00192281e6c555fd0;
	//wire [511:0] data = 512'h0;
	//wire [511:0] data = {256'h0000010000000000000000000000000000000000000000000000000080000000, 256'h0};
	//wire [255:0] data = 256'h0;
	//wire [0:511] data = 512'hc13858e5a13de1500e54a1c85f0132e688e131b93d7bf9a00192281e6c555fd0c13858e5a13de1500e54a1c85f0132e688e131b93d7bf9a00192281e6c555fd0;
	//wire [511:0] data = 512'h00000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000100;
	//wire [511:0] data = 512'hDEADBEEF000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000100;
	wire [511:0] data =   512'hdeadbeefcafe00000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000170;

	wire [511:0] data_end_rev;
	//assign data_rev = data;
	wire [255:0] hash_out;
	genvar i;
	generate
		for (i=0; i<16; i=i+1) begin: ENDIAN_REV
			assign data_end_rev[32*i +: 32] = data[32*(15-i) +: 32];
		end
	endgenerate
	//   00000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000100;
	//	5be0cd191f83d9ab9b05688c510e527fa54ff53a3c6ef372bb67ae856a09e667
	
	always 
	begin
		#5 clk = ~clk;
	end

//6a09e667bb67ae853c6ef372a54ff53a510e527f9b05688c1f83d9ab5be0cd19

//5be0cd191f83d9ab9b05688c510e527fa54ff53a3c6ef372bb67ae856a09e667

	sha256_transform #(.LOOP(LOOP)) uut (
		.clk(clk),
		.feedback(1'b0),
		.cnt(6'd0),
		//.rx_state(256'h6a09e667bb67ae853c6ef372a54ff53a510e527f9b05688c1f83d9ab5be0cd19),
		.rx_state(256'h5be0cd191f83d9ab9b05688c510e527fa54ff53a3c6ef372bb67ae856a09e667),
		//.rx_input(data),
		.rx_input(data_end_rev),
		//.rx_input({256'h0000010000000000000000000000000000000000000000000000000080000000, data}),
		//.rx_input({256'h00000000000000000000000000000000800000000000000000000000000000010
		//.rx_input({256'h80000000000000000000000000000000000000000000000000000000000000020, data}),
		.tx_hash(hash_out)
	);

	wire [255:0] hash_out_rev;
	generate
		for (i=0; i<8; i=i+1) begin: HASH_OUT_REV
			assign hash_out_rev[32*i +: 32] = hash_out[32*(7-i) +: 32];
		end
	endgenerate

	always@(posedge clk)
	begin
		$display("hashinp=%x", data);
		$display("hashirev=%x", data_end_rev);
		$display("hashout=%x", hash_out);
		$display("hashorev=%x", hash_out_rev);
	end
endmodule
